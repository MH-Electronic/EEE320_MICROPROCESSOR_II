// MicroP.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module MicroP (
		input  wire       bluetooth_uart_rxd,    // bluetooth_uart.rxd
		output wire       bluetooth_uart_txd,    //               .txd
		input  wire       button_int_export,     //     button_int.export
		output wire       buzzer_export,         //         buzzer.export
		input  wire       clk_clk,               //            clk.clk
		output wire       clk_25_export,         //         clk_25.export
		output wire       clk_check_export,      //      clk_check.export
		input  wire [3:0] keypad_column_export,  //  keypad_column.export
		output wire [3:0] keypad_row_export,     //     keypad_row.export
		input  wire       reset_reset_n,         //          reset.reset_n
		output wire       rfid_cs_export,        //        rfid_cs.export
		input  wire       rfid_spi_MISO,         //       rfid_spi.MISO
		output wire       rfid_spi_MOSI,         //               .MOSI
		output wire       rfid_spi_SCLK,         //               .SCLK
		output wire       rfid_spi_SS_n,         //               .SS_n
		input  wire [7:0] switches_export,       //       switches.export
		input  wire       ultrasonic_in_export,  //  ultrasonic_in.export
		output wire       ultrasonic_out_export, // ultrasonic_out.export
		output wire       vga_external_CLK,      //   vga_external.CLK
		output wire       vga_external_HS,       //               .HS
		output wire       vga_external_VS,       //               .VS
		output wire       vga_external_BLANK,    //               .BLANK
		output wire       vga_external_SYNC,     //               .SYNC
		output wire [7:0] vga_external_R,        //               .R
		output wire [7:0] vga_external_G,        //               .G
		output wire [7:0] vga_external_B         //               .B
	);

	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                               // video_character_buffer_with_dma_0:stream_valid -> vga_controller:valid
	wire  [29:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                // video_character_buffer_with_dma_0:stream_data -> vga_controller:data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                               // vga_controller:ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                       // video_character_buffer_with_dma_0:stream_startofpacket -> vga_controller:startofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                         // video_character_buffer_with_dma_0:stream_endofpacket -> vga_controller:endofpacket
	wire         clk_25_outclk0_clk;                                                                       // clk_25:outclk_0 -> [mm_interconnect_0:clk_25_outclk0_clk, rst_controller_002:clk, vga_controller:clk, video_character_buffer_with_dma_0:clk]
	wire  [31:0] nios2_data_master_readdata;                                                               // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                                            // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                                            // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [16:0] nios2_data_master_address;                                                                // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                                             // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                                   // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                                                  // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                                              // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                                        // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                                     // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [16:0] nios2_instruction_master_address;                                                         // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                                            // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;    // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest; // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;   // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;    // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;      // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                                      // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                                        // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                                     // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                                         // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                            // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                                           // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                                       // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                                      // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                                       // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                                         // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                                      // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                                      // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                                          // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                                             // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                                       // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                                            // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                                        // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_clk_check_s1_chipselect;                                                // mm_interconnect_0:Clk_check_s1_chipselect -> Clk_check:chipselect
	wire  [31:0] mm_interconnect_0_clk_check_s1_readdata;                                                  // Clk_check:readdata -> mm_interconnect_0:Clk_check_s1_readdata
	wire   [1:0] mm_interconnect_0_clk_check_s1_address;                                                   // mm_interconnect_0:Clk_check_s1_address -> Clk_check:address
	wire         mm_interconnect_0_clk_check_s1_write;                                                     // mm_interconnect_0:Clk_check_s1_write -> Clk_check:write_n
	wire  [31:0] mm_interconnect_0_clk_check_s1_writedata;                                                 // mm_interconnect_0:Clk_check_s1_writedata -> Clk_check:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                                                   // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                                                    // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire         mm_interconnect_0_ram_s1_chipselect;                                                      // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                                        // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [13:0] mm_interconnect_0_ram_s1_address;                                                         // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                                                      // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                                           // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                                       // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                                           // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_bluetooth_uart_s1_chipselect;                                           // mm_interconnect_0:bluetooth_UART_s1_chipselect -> bluetooth_UART:chipselect
	wire  [15:0] mm_interconnect_0_bluetooth_uart_s1_readdata;                                             // bluetooth_UART:readdata -> mm_interconnect_0:bluetooth_UART_s1_readdata
	wire   [2:0] mm_interconnect_0_bluetooth_uart_s1_address;                                              // mm_interconnect_0:bluetooth_UART_s1_address -> bluetooth_UART:address
	wire         mm_interconnect_0_bluetooth_uart_s1_read;                                                 // mm_interconnect_0:bluetooth_UART_s1_read -> bluetooth_UART:read_n
	wire         mm_interconnect_0_bluetooth_uart_s1_begintransfer;                                        // mm_interconnect_0:bluetooth_UART_s1_begintransfer -> bluetooth_UART:begintransfer
	wire         mm_interconnect_0_bluetooth_uart_s1_write;                                                // mm_interconnect_0:bluetooth_UART_s1_write -> bluetooth_UART:write_n
	wire  [15:0] mm_interconnect_0_bluetooth_uart_s1_writedata;                                            // mm_interconnect_0:bluetooth_UART_s1_writedata -> bluetooth_UART:writedata
	wire  [31:0] mm_interconnect_0_keypad_column_s1_readdata;                                              // keypad_column:readdata -> mm_interconnect_0:keypad_column_s1_readdata
	wire   [1:0] mm_interconnect_0_keypad_column_s1_address;                                               // mm_interconnect_0:keypad_column_s1_address -> keypad_column:address
	wire         mm_interconnect_0_button_int_s1_chipselect;                                               // mm_interconnect_0:button_int_s1_chipselect -> button_int:chipselect
	wire  [31:0] mm_interconnect_0_button_int_s1_readdata;                                                 // button_int:readdata -> mm_interconnect_0:button_int_s1_readdata
	wire   [1:0] mm_interconnect_0_button_int_s1_address;                                                  // mm_interconnect_0:button_int_s1_address -> button_int:address
	wire         mm_interconnect_0_button_int_s1_write;                                                    // mm_interconnect_0:button_int_s1_write -> button_int:write_n
	wire  [31:0] mm_interconnect_0_button_int_s1_writedata;                                                // mm_interconnect_0:button_int_s1_writedata -> button_int:writedata
	wire         mm_interconnect_0_buzzer_s1_chipselect;                                                   // mm_interconnect_0:Buzzer_s1_chipselect -> Buzzer:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                                                     // Buzzer:readdata -> mm_interconnect_0:Buzzer_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                                                      // mm_interconnect_0:Buzzer_s1_address -> Buzzer:address
	wire         mm_interconnect_0_buzzer_s1_write;                                                        // mm_interconnect_0:Buzzer_s1_write -> Buzzer:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                                                    // mm_interconnect_0:Buzzer_s1_writedata -> Buzzer:writedata
	wire         mm_interconnect_0_ultrasonic_out_s1_chipselect;                                           // mm_interconnect_0:ultrasonic_out_s1_chipselect -> ultrasonic_out:chipselect
	wire  [31:0] mm_interconnect_0_ultrasonic_out_s1_readdata;                                             // ultrasonic_out:readdata -> mm_interconnect_0:ultrasonic_out_s1_readdata
	wire   [1:0] mm_interconnect_0_ultrasonic_out_s1_address;                                              // mm_interconnect_0:ultrasonic_out_s1_address -> ultrasonic_out:address
	wire         mm_interconnect_0_ultrasonic_out_s1_write;                                                // mm_interconnect_0:ultrasonic_out_s1_write -> ultrasonic_out:write_n
	wire  [31:0] mm_interconnect_0_ultrasonic_out_s1_writedata;                                            // mm_interconnect_0:ultrasonic_out_s1_writedata -> ultrasonic_out:writedata
	wire         mm_interconnect_0_keypad_row_s1_chipselect;                                               // mm_interconnect_0:keypad_row_s1_chipselect -> keypad_row:chipselect
	wire  [31:0] mm_interconnect_0_keypad_row_s1_readdata;                                                 // keypad_row:readdata -> mm_interconnect_0:keypad_row_s1_readdata
	wire   [1:0] mm_interconnect_0_keypad_row_s1_address;                                                  // mm_interconnect_0:keypad_row_s1_address -> keypad_row:address
	wire         mm_interconnect_0_keypad_row_s1_write;                                                    // mm_interconnect_0:keypad_row_s1_write -> keypad_row:write_n
	wire  [31:0] mm_interconnect_0_keypad_row_s1_writedata;                                                // mm_interconnect_0:keypad_row_s1_writedata -> keypad_row:writedata
	wire         mm_interconnect_0_rfid_cs_s1_chipselect;                                                  // mm_interconnect_0:RFID_cs_s1_chipselect -> RFID_cs:chipselect
	wire  [31:0] mm_interconnect_0_rfid_cs_s1_readdata;                                                    // RFID_cs:readdata -> mm_interconnect_0:RFID_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_rfid_cs_s1_address;                                                     // mm_interconnect_0:RFID_cs_s1_address -> RFID_cs:address
	wire         mm_interconnect_0_rfid_cs_s1_write;                                                       // mm_interconnect_0:RFID_cs_s1_write -> RFID_cs:write_n
	wire  [31:0] mm_interconnect_0_rfid_cs_s1_writedata;                                                   // mm_interconnect_0:RFID_cs_s1_writedata -> RFID_cs:writedata
	wire  [31:0] mm_interconnect_0_ultrasonic_in_s1_readdata;                                              // ultrasonic_in:readdata -> mm_interconnect_0:ultrasonic_in_s1_readdata
	wire   [1:0] mm_interconnect_0_ultrasonic_in_s1_address;                                               // mm_interconnect_0:ultrasonic_in_s1_address -> ultrasonic_in:address
	wire         mm_interconnect_0_rfid_spi_spi_control_port_chipselect;                                   // mm_interconnect_0:RFID_spi_spi_control_port_chipselect -> RFID_spi:spi_select
	wire  [15:0] mm_interconnect_0_rfid_spi_spi_control_port_readdata;                                     // RFID_spi:data_to_cpu -> mm_interconnect_0:RFID_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_rfid_spi_spi_control_port_address;                                      // mm_interconnect_0:RFID_spi_spi_control_port_address -> RFID_spi:mem_addr
	wire         mm_interconnect_0_rfid_spi_spi_control_port_read;                                         // mm_interconnect_0:RFID_spi_spi_control_port_read -> RFID_spi:read_n
	wire         mm_interconnect_0_rfid_spi_spi_control_port_write;                                        // mm_interconnect_0:RFID_spi_spi_control_port_write -> RFID_spi:write_n
	wire  [15:0] mm_interconnect_0_rfid_spi_spi_control_port_writedata;                                    // mm_interconnect_0:RFID_spi_spi_control_port_writedata -> RFID_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                                 // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                 // bluetooth_UART:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                 // button_int:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                 // RFID_spi:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_irq_irq;                                                                            // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [Buzzer:reset_n, bluetooth_UART:reset_n, mm_interconnect_0:sysid_qsys_reset_reset_bridge_in_reset_reset, sysid_qsys:reset_n]
	wire         rst_controller_001_reset_out_reset;                                                       // rst_controller_001:reset_out -> [Clk_check:reset_n, RFID_cs:reset_n, RFID_spi:reset_n, Switches:reset_n, button_int:reset_n, irq_mapper:reset, jtag:rst_n, keypad_column:reset_n, keypad_row:reset_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, ram:reset, rst_translator:in_reset, ultrasonic_in:reset_n, ultrasonic_out:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                                   // rst_controller_001:reset_req -> [nios2:reset_req, ram:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                                                          // nios2:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                                                       // rst_controller_002:reset_out -> [mm_interconnect_0:video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset, vga_controller:reset, video_character_buffer_with_dma_0:reset]

	MicroP_Buzzer buzzer (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                           // external_connection.export
	);

	MicroP_Buzzer clk_check (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_clk_check_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clk_check_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clk_check_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clk_check_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clk_check_s1_readdata),   //                    .readdata
		.out_port   (clk_check_export)                           // external_connection.export
	);

	MicroP_Buzzer rfid_cs (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_rfid_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rfid_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rfid_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rfid_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rfid_cs_s1_readdata),   //                    .readdata
		.out_port   (rfid_cs_export)                           // external_connection.export
	);

	MicroP_RFID_spi rfid_spi (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_rfid_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_rfid_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_rfid_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_rfid_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_rfid_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_rfid_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                               //              irq.irq
		.MISO          (rfid_spi_MISO),                                          //         external.export
		.MOSI          (rfid_spi_MOSI),                                          //                 .export
		.SCLK          (rfid_spi_SCLK),                                          //                 .export
		.SS_n          (rfid_spi_SS_n)                                           //                 .export
	);

	MicroP_Switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	MicroP_bluetooth_UART bluetooth_uart (
		.clk           (clk_clk),                                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address       (mm_interconnect_0_bluetooth_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_bluetooth_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_bluetooth_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_bluetooth_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_bluetooth_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_bluetooth_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_bluetooth_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                                  //                    .dataavailable
		.readyfordata  (),                                                  //                    .readyfordata
		.rxd           (bluetooth_uart_rxd),                                // external_connection.export
		.txd           (bluetooth_uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver1_irq)                           //                 irq.irq
	);

	MicroP_button_int button_int (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_int_s1_readdata),   //                    .readdata
		.in_port    (button_int_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	MicroP_clk_25 clk_25 (
		.refclk   (clk_clk),            //  refclk.clk
		.rst      (~reset_reset_n),     //   reset.reset
		.outclk_0 (clk_25_outclk0_clk), // outclk0.clk
		.locked   (clk_25_export)       //  locked.export
	);

	MicroP_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	MicroP_keypad_column keypad_column (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_keypad_column_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keypad_column_s1_readdata), //                    .readdata
		.in_port  (keypad_column_export)                         // external_connection.export
	);

	MicroP_keypad_row keypad_row (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_keypad_row_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keypad_row_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keypad_row_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keypad_row_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keypad_row_s1_readdata),   //                    .readdata
		.out_port   (keypad_row_export)                           // external_connection.export
	);

	MicroP_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	MicroP_ram ram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),         //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)  //       .reset_req
	);

	MicroP_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	MicroP_ultrasonic_in ultrasonic_in (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_ultrasonic_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ultrasonic_in_s1_readdata), //                    .readdata
		.in_port  (ultrasonic_in_export)                         // external_connection.export
	);

	MicroP_Buzzer ultrasonic_out (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_ultrasonic_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ultrasonic_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ultrasonic_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ultrasonic_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ultrasonic_out_s1_readdata),   //                    .readdata
		.out_port   (ultrasonic_out_export)                           // external_connection.export
	);

	MicroP_vga_controller vga_controller (
		.clk           (clk_25_outclk0_clk),                                                 //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                                 //              reset.reset
		.data          (video_character_buffer_with_dma_0_avalon_char_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                   .endofpacket
		.valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                   .valid
		.ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                   .ready
		.VGA_CLK       (vga_external_CLK),                                                   // external_interface.export
		.VGA_HS        (vga_external_HS),                                                    //                   .export
		.VGA_VS        (vga_external_VS),                                                    //                   .export
		.VGA_BLANK     (vga_external_BLANK),                                                 //                   .export
		.VGA_SYNC      (vga_external_SYNC),                                                  //                   .export
		.VGA_R         (vga_external_R),                                                     //                   .export
		.VGA_G         (vga_external_G),                                                     //                   .export
		.VGA_B         (vga_external_B)                                                      //                   .export
	);

	MicroP_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clk_25_outclk0_clk),                                                                       //                       clk.clk
		.reset                (rst_controller_002_reset_out_reset),                                                       //                     reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	MicroP_mm_interconnect_0 mm_interconnect_0 (
		.clk_25_outclk0_clk                                                     (clk_25_outclk0_clk),                                                                       //                                                clk_25_outclk0.clk
		.system_clk_clk_clk                                                     (clk_clk),                                                                                  //                                                system_clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset                                (rst_controller_001_reset_out_reset),                                                       //                             nios2_reset_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset                           (rst_controller_reset_out_reset),                                                           //                        sysid_qsys_reset_reset_bridge_in_reset.reset
		.video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                                                       // video_character_buffer_with_dma_0_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                                              (nios2_data_master_address),                                                                //                                             nios2_data_master.address
		.nios2_data_master_waitrequest                                          (nios2_data_master_waitrequest),                                                            //                                                              .waitrequest
		.nios2_data_master_byteenable                                           (nios2_data_master_byteenable),                                                             //                                                              .byteenable
		.nios2_data_master_read                                                 (nios2_data_master_read),                                                                   //                                                              .read
		.nios2_data_master_readdata                                             (nios2_data_master_readdata),                                                               //                                                              .readdata
		.nios2_data_master_write                                                (nios2_data_master_write),                                                                  //                                                              .write
		.nios2_data_master_writedata                                            (nios2_data_master_writedata),                                                              //                                                              .writedata
		.nios2_data_master_debugaccess                                          (nios2_data_master_debugaccess),                                                            //                                                              .debugaccess
		.nios2_instruction_master_address                                       (nios2_instruction_master_address),                                                         //                                      nios2_instruction_master.address
		.nios2_instruction_master_waitrequest                                   (nios2_instruction_master_waitrequest),                                                     //                                                              .waitrequest
		.nios2_instruction_master_read                                          (nios2_instruction_master_read),                                                            //                                                              .read
		.nios2_instruction_master_readdata                                      (nios2_instruction_master_readdata),                                                        //                                                              .readdata
		.bluetooth_UART_s1_address                                              (mm_interconnect_0_bluetooth_uart_s1_address),                                              //                                             bluetooth_UART_s1.address
		.bluetooth_UART_s1_write                                                (mm_interconnect_0_bluetooth_uart_s1_write),                                                //                                                              .write
		.bluetooth_UART_s1_read                                                 (mm_interconnect_0_bluetooth_uart_s1_read),                                                 //                                                              .read
		.bluetooth_UART_s1_readdata                                             (mm_interconnect_0_bluetooth_uart_s1_readdata),                                             //                                                              .readdata
		.bluetooth_UART_s1_writedata                                            (mm_interconnect_0_bluetooth_uart_s1_writedata),                                            //                                                              .writedata
		.bluetooth_UART_s1_begintransfer                                        (mm_interconnect_0_bluetooth_uart_s1_begintransfer),                                        //                                                              .begintransfer
		.bluetooth_UART_s1_chipselect                                           (mm_interconnect_0_bluetooth_uart_s1_chipselect),                                           //                                                              .chipselect
		.button_int_s1_address                                                  (mm_interconnect_0_button_int_s1_address),                                                  //                                                 button_int_s1.address
		.button_int_s1_write                                                    (mm_interconnect_0_button_int_s1_write),                                                    //                                                              .write
		.button_int_s1_readdata                                                 (mm_interconnect_0_button_int_s1_readdata),                                                 //                                                              .readdata
		.button_int_s1_writedata                                                (mm_interconnect_0_button_int_s1_writedata),                                                //                                                              .writedata
		.button_int_s1_chipselect                                               (mm_interconnect_0_button_int_s1_chipselect),                                               //                                                              .chipselect
		.Buzzer_s1_address                                                      (mm_interconnect_0_buzzer_s1_address),                                                      //                                                     Buzzer_s1.address
		.Buzzer_s1_write                                                        (mm_interconnect_0_buzzer_s1_write),                                                        //                                                              .write
		.Buzzer_s1_readdata                                                     (mm_interconnect_0_buzzer_s1_readdata),                                                     //                                                              .readdata
		.Buzzer_s1_writedata                                                    (mm_interconnect_0_buzzer_s1_writedata),                                                    //                                                              .writedata
		.Buzzer_s1_chipselect                                                   (mm_interconnect_0_buzzer_s1_chipselect),                                                   //                                                              .chipselect
		.Clk_check_s1_address                                                   (mm_interconnect_0_clk_check_s1_address),                                                   //                                                  Clk_check_s1.address
		.Clk_check_s1_write                                                     (mm_interconnect_0_clk_check_s1_write),                                                     //                                                              .write
		.Clk_check_s1_readdata                                                  (mm_interconnect_0_clk_check_s1_readdata),                                                  //                                                              .readdata
		.Clk_check_s1_writedata                                                 (mm_interconnect_0_clk_check_s1_writedata),                                                 //                                                              .writedata
		.Clk_check_s1_chipselect                                                (mm_interconnect_0_clk_check_s1_chipselect),                                                //                                                              .chipselect
		.jtag_avalon_jtag_slave_address                                         (mm_interconnect_0_jtag_avalon_jtag_slave_address),                                         //                                        jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                                           (mm_interconnect_0_jtag_avalon_jtag_slave_write),                                           //                                                              .write
		.jtag_avalon_jtag_slave_read                                            (mm_interconnect_0_jtag_avalon_jtag_slave_read),                                            //                                                              .read
		.jtag_avalon_jtag_slave_readdata                                        (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                                        //                                                              .readdata
		.jtag_avalon_jtag_slave_writedata                                       (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                                       //                                                              .writedata
		.jtag_avalon_jtag_slave_waitrequest                                     (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                                     //                                                              .waitrequest
		.jtag_avalon_jtag_slave_chipselect                                      (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                                      //                                                              .chipselect
		.keypad_column_s1_address                                               (mm_interconnect_0_keypad_column_s1_address),                                               //                                              keypad_column_s1.address
		.keypad_column_s1_readdata                                              (mm_interconnect_0_keypad_column_s1_readdata),                                              //                                                              .readdata
		.keypad_row_s1_address                                                  (mm_interconnect_0_keypad_row_s1_address),                                                  //                                                 keypad_row_s1.address
		.keypad_row_s1_write                                                    (mm_interconnect_0_keypad_row_s1_write),                                                    //                                                              .write
		.keypad_row_s1_readdata                                                 (mm_interconnect_0_keypad_row_s1_readdata),                                                 //                                                              .readdata
		.keypad_row_s1_writedata                                                (mm_interconnect_0_keypad_row_s1_writedata),                                                //                                                              .writedata
		.keypad_row_s1_chipselect                                               (mm_interconnect_0_keypad_row_s1_chipselect),                                               //                                                              .chipselect
		.nios2_debug_mem_slave_address                                          (mm_interconnect_0_nios2_debug_mem_slave_address),                                          //                                         nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                                            (mm_interconnect_0_nios2_debug_mem_slave_write),                                            //                                                              .write
		.nios2_debug_mem_slave_read                                             (mm_interconnect_0_nios2_debug_mem_slave_read),                                             //                                                              .read
		.nios2_debug_mem_slave_readdata                                         (mm_interconnect_0_nios2_debug_mem_slave_readdata),                                         //                                                              .readdata
		.nios2_debug_mem_slave_writedata                                        (mm_interconnect_0_nios2_debug_mem_slave_writedata),                                        //                                                              .writedata
		.nios2_debug_mem_slave_byteenable                                       (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                                       //                                                              .byteenable
		.nios2_debug_mem_slave_waitrequest                                      (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                                      //                                                              .waitrequest
		.nios2_debug_mem_slave_debugaccess                                      (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                                      //                                                              .debugaccess
		.ram_s1_address                                                         (mm_interconnect_0_ram_s1_address),                                                         //                                                        ram_s1.address
		.ram_s1_write                                                           (mm_interconnect_0_ram_s1_write),                                                           //                                                              .write
		.ram_s1_readdata                                                        (mm_interconnect_0_ram_s1_readdata),                                                        //                                                              .readdata
		.ram_s1_writedata                                                       (mm_interconnect_0_ram_s1_writedata),                                                       //                                                              .writedata
		.ram_s1_byteenable                                                      (mm_interconnect_0_ram_s1_byteenable),                                                      //                                                              .byteenable
		.ram_s1_chipselect                                                      (mm_interconnect_0_ram_s1_chipselect),                                                      //                                                              .chipselect
		.ram_s1_clken                                                           (mm_interconnect_0_ram_s1_clken),                                                           //                                                              .clken
		.RFID_cs_s1_address                                                     (mm_interconnect_0_rfid_cs_s1_address),                                                     //                                                    RFID_cs_s1.address
		.RFID_cs_s1_write                                                       (mm_interconnect_0_rfid_cs_s1_write),                                                       //                                                              .write
		.RFID_cs_s1_readdata                                                    (mm_interconnect_0_rfid_cs_s1_readdata),                                                    //                                                              .readdata
		.RFID_cs_s1_writedata                                                   (mm_interconnect_0_rfid_cs_s1_writedata),                                                   //                                                              .writedata
		.RFID_cs_s1_chipselect                                                  (mm_interconnect_0_rfid_cs_s1_chipselect),                                                  //                                                              .chipselect
		.RFID_spi_spi_control_port_address                                      (mm_interconnect_0_rfid_spi_spi_control_port_address),                                      //                                     RFID_spi_spi_control_port.address
		.RFID_spi_spi_control_port_write                                        (mm_interconnect_0_rfid_spi_spi_control_port_write),                                        //                                                              .write
		.RFID_spi_spi_control_port_read                                         (mm_interconnect_0_rfid_spi_spi_control_port_read),                                         //                                                              .read
		.RFID_spi_spi_control_port_readdata                                     (mm_interconnect_0_rfid_spi_spi_control_port_readdata),                                     //                                                              .readdata
		.RFID_spi_spi_control_port_writedata                                    (mm_interconnect_0_rfid_spi_spi_control_port_writedata),                                    //                                                              .writedata
		.RFID_spi_spi_control_port_chipselect                                   (mm_interconnect_0_rfid_spi_spi_control_port_chipselect),                                   //                                                              .chipselect
		.Switches_s1_address                                                    (mm_interconnect_0_switches_s1_address),                                                    //                                                   Switches_s1.address
		.Switches_s1_readdata                                                   (mm_interconnect_0_switches_s1_readdata),                                                   //                                                              .readdata
		.sysid_qsys_control_slave_address                                       (mm_interconnect_0_sysid_qsys_control_slave_address),                                       //                                      sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                      (mm_interconnect_0_sysid_qsys_control_slave_readdata),                                      //                                                              .readdata
		.ultrasonic_in_s1_address                                               (mm_interconnect_0_ultrasonic_in_s1_address),                                               //                                              ultrasonic_in_s1.address
		.ultrasonic_in_s1_readdata                                              (mm_interconnect_0_ultrasonic_in_s1_readdata),                                              //                                                              .readdata
		.ultrasonic_out_s1_address                                              (mm_interconnect_0_ultrasonic_out_s1_address),                                              //                                             ultrasonic_out_s1.address
		.ultrasonic_out_s1_write                                                (mm_interconnect_0_ultrasonic_out_s1_write),                                                //                                                              .write
		.ultrasonic_out_s1_readdata                                             (mm_interconnect_0_ultrasonic_out_s1_readdata),                                             //                                                              .readdata
		.ultrasonic_out_s1_writedata                                            (mm_interconnect_0_ultrasonic_out_s1_writedata),                                            //                                                              .writedata
		.ultrasonic_out_s1_chipselect                                           (mm_interconnect_0_ultrasonic_out_s1_chipselect),                                           //                                                              .chipselect
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //    video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                                                              .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                                                              .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                                                              .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                                                              .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //                                                              .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                                                              .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                                                              .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    //   video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                                                              .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                                                              .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                                                              .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                                                              .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                                                              .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect)  //                                                              .chipselect
	);

	MicroP_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),        // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_25_outclk0_clk),                 //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
